`timescale 1ns / 1ns

module cpu_pc(
    input               clock,
    input               reset,
    input               stall,
    input               p2_pipeline_bubble,

    // Connection to execution unit
    input               p3_jump,
    input [31:0]        p3_jump_target,

    // Connection to instruction bus
    output reg [31:0]   p1_pc,
    output reg [31:0]   p2_pc,
    output reg [31:0]   p3_pc
);

always @(*) begin
    if (p3_jump)
        p1_pc = p3_jump_target;
    else if (p2_pipeline_bubble || stall)
        p1_pc = p2_pc;
    else
        p1_pc = p2_pc + 4;

    if (reset) begin
        p1_pc = 32'hffff0000;
    end
end


always @(posedge clock) begin
    if (!stall) begin
        p2_pc <= p1_pc;
        p3_pc <= p2_pc;
    end
end

// synthesis translate_off
always @(posedge clock) begin
    if (p2_pc == 32'h0) begin
        @(posedge clock);
        $finish();
    end
end
// synthesis translate_on


endmodule